module tt_um_roy1707018_ro2 (clk,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uo_out);
 input clk;
 input rst_n;
 input VPWR;
 input VGND;
 input [7:0] ui_in;
 output [7:0] uo_out;

 wire _00_;
 wire _01_;
 wire \u_ro_only.ro_gen[0].ro1.cq4 ;
 wire \u_ro_only.ro_gen[0].ro1.en ;
 wire \u_ro_only.ro_gen[0].ro1.q ;
 wire \u_ro_only.ro_gen[0].ro1.q0 ;
 wire \u_ro_only.ro_gen[0].ro1.q1 ;
 wire \u_ro_only.ro_gen[0].ro1.q2 ;
 wire \u_ro_only.ro_gen[0].ro1.q3 ;
 wire \u_ro_only.ro_gen[0].ro1.q4 ;
 wire \u_ro_only.ro_gen[0].ro2.cq4 ;
 wire \u_ro_only.ro_gen[0].ro2.en ;
 wire \u_ro_only.ro_gen[0].ro2.q ;
 wire \u_ro_only.ro_gen[0].ro2.q0 ;
 wire \u_ro_only.ro_gen[0].ro2.q1 ;
 wire \u_ro_only.ro_gen[0].ro2.q2 ;
 wire \u_ro_only.ro_gen[0].ro2.q3 ;
 wire \u_ro_only.ro_gen[0].ro2.q4 ;
 wire \u_ro_only.ro_gen[10].ro1.cq4 ;
 wire \u_ro_only.ro_gen[10].ro1.q ;
 wire \u_ro_only.ro_gen[10].ro1.q0 ;
 wire \u_ro_only.ro_gen[10].ro1.q1 ;
 wire \u_ro_only.ro_gen[10].ro1.q2 ;
 wire \u_ro_only.ro_gen[10].ro1.q3 ;
 wire \u_ro_only.ro_gen[10].ro1.q4 ;
 wire \u_ro_only.ro_gen[10].ro2.cq4 ;
 wire \u_ro_only.ro_gen[10].ro2.q ;
 wire \u_ro_only.ro_gen[10].ro2.q0 ;
 wire \u_ro_only.ro_gen[10].ro2.q1 ;
 wire \u_ro_only.ro_gen[10].ro2.q2 ;
 wire \u_ro_only.ro_gen[10].ro2.q3 ;
 wire \u_ro_only.ro_gen[10].ro2.q4 ;
 wire \u_ro_only.ro_gen[11].ro1.cq4 ;
 wire \u_ro_only.ro_gen[11].ro1.q ;
 wire \u_ro_only.ro_gen[11].ro1.q0 ;
 wire \u_ro_only.ro_gen[11].ro1.q1 ;
 wire \u_ro_only.ro_gen[11].ro1.q2 ;
 wire \u_ro_only.ro_gen[11].ro1.q3 ;
 wire \u_ro_only.ro_gen[11].ro1.q4 ;
 wire \u_ro_only.ro_gen[11].ro2.cq4 ;
 wire \u_ro_only.ro_gen[11].ro2.q ;
 wire \u_ro_only.ro_gen[11].ro2.q0 ;
 wire \u_ro_only.ro_gen[11].ro2.q1 ;
 wire \u_ro_only.ro_gen[11].ro2.q2 ;
 wire \u_ro_only.ro_gen[11].ro2.q3 ;
 wire \u_ro_only.ro_gen[11].ro2.q4 ;
 wire \u_ro_only.ro_gen[12].ro1.cq4 ;
 wire \u_ro_only.ro_gen[12].ro1.q ;
 wire \u_ro_only.ro_gen[12].ro1.q0 ;
 wire \u_ro_only.ro_gen[12].ro1.q1 ;
 wire \u_ro_only.ro_gen[12].ro1.q2 ;
 wire \u_ro_only.ro_gen[12].ro1.q3 ;
 wire \u_ro_only.ro_gen[12].ro1.q4 ;
 wire \u_ro_only.ro_gen[12].ro2.cq4 ;
 wire \u_ro_only.ro_gen[12].ro2.q ;
 wire \u_ro_only.ro_gen[12].ro2.q0 ;
 wire \u_ro_only.ro_gen[12].ro2.q1 ;
 wire \u_ro_only.ro_gen[12].ro2.q2 ;
 wire \u_ro_only.ro_gen[12].ro2.q3 ;
 wire \u_ro_only.ro_gen[12].ro2.q4 ;
 wire \u_ro_only.ro_gen[13].ro1.cq4 ;
 wire \u_ro_only.ro_gen[13].ro1.q ;
 wire \u_ro_only.ro_gen[13].ro1.q0 ;
 wire \u_ro_only.ro_gen[13].ro1.q1 ;
 wire \u_ro_only.ro_gen[13].ro1.q2 ;
 wire \u_ro_only.ro_gen[13].ro1.q3 ;
 wire \u_ro_only.ro_gen[13].ro1.q4 ;
 wire \u_ro_only.ro_gen[13].ro2.cq4 ;
 wire \u_ro_only.ro_gen[13].ro2.q ;
 wire \u_ro_only.ro_gen[13].ro2.q0 ;
 wire \u_ro_only.ro_gen[13].ro2.q1 ;
 wire \u_ro_only.ro_gen[13].ro2.q2 ;
 wire \u_ro_only.ro_gen[13].ro2.q3 ;
 wire \u_ro_only.ro_gen[13].ro2.q4 ;
 wire \u_ro_only.ro_gen[14].ro1.cq4 ;
 wire \u_ro_only.ro_gen[14].ro1.q ;
 wire \u_ro_only.ro_gen[14].ro1.q0 ;
 wire \u_ro_only.ro_gen[14].ro1.q1 ;
 wire \u_ro_only.ro_gen[14].ro1.q2 ;
 wire \u_ro_only.ro_gen[14].ro1.q3 ;
 wire \u_ro_only.ro_gen[14].ro1.q4 ;
 wire \u_ro_only.ro_gen[14].ro2.cq4 ;
 wire \u_ro_only.ro_gen[14].ro2.q ;
 wire \u_ro_only.ro_gen[14].ro2.q0 ;
 wire \u_ro_only.ro_gen[14].ro2.q1 ;
 wire \u_ro_only.ro_gen[14].ro2.q2 ;
 wire \u_ro_only.ro_gen[14].ro2.q3 ;
 wire \u_ro_only.ro_gen[14].ro2.q4 ;
 wire \u_ro_only.ro_gen[15].ro1.cq4 ;
 wire \u_ro_only.ro_gen[15].ro1.q ;
 wire \u_ro_only.ro_gen[15].ro1.q0 ;
 wire \u_ro_only.ro_gen[15].ro1.q1 ;
 wire \u_ro_only.ro_gen[15].ro1.q2 ;
 wire \u_ro_only.ro_gen[15].ro1.q3 ;
 wire \u_ro_only.ro_gen[15].ro1.q4 ;
 wire \u_ro_only.ro_gen[15].ro2.cq4 ;
 wire \u_ro_only.ro_gen[15].ro2.q ;
 wire \u_ro_only.ro_gen[15].ro2.q0 ;
 wire \u_ro_only.ro_gen[15].ro2.q1 ;
 wire \u_ro_only.ro_gen[15].ro2.q2 ;
 wire \u_ro_only.ro_gen[15].ro2.q3 ;
 wire \u_ro_only.ro_gen[15].ro2.q4 ;
 wire \u_ro_only.ro_gen[1].ro1.cq4 ;
 wire \u_ro_only.ro_gen[1].ro1.q ;
 wire \u_ro_only.ro_gen[1].ro1.q0 ;
 wire \u_ro_only.ro_gen[1].ro1.q1 ;
 wire \u_ro_only.ro_gen[1].ro1.q2 ;
 wire \u_ro_only.ro_gen[1].ro1.q3 ;
 wire \u_ro_only.ro_gen[1].ro1.q4 ;
 wire \u_ro_only.ro_gen[1].ro2.cq4 ;
 wire \u_ro_only.ro_gen[1].ro2.q ;
 wire \u_ro_only.ro_gen[1].ro2.q0 ;
 wire \u_ro_only.ro_gen[1].ro2.q1 ;
 wire \u_ro_only.ro_gen[1].ro2.q2 ;
 wire \u_ro_only.ro_gen[1].ro2.q3 ;
 wire \u_ro_only.ro_gen[1].ro2.q4 ;
 wire \u_ro_only.ro_gen[2].ro1.cq4 ;
 wire \u_ro_only.ro_gen[2].ro1.q ;
 wire \u_ro_only.ro_gen[2].ro1.q0 ;
 wire \u_ro_only.ro_gen[2].ro1.q1 ;
 wire \u_ro_only.ro_gen[2].ro1.q2 ;
 wire \u_ro_only.ro_gen[2].ro1.q3 ;
 wire \u_ro_only.ro_gen[2].ro1.q4 ;
 wire \u_ro_only.ro_gen[2].ro2.cq4 ;
 wire \u_ro_only.ro_gen[2].ro2.q ;
 wire \u_ro_only.ro_gen[2].ro2.q0 ;
 wire \u_ro_only.ro_gen[2].ro2.q1 ;
 wire \u_ro_only.ro_gen[2].ro2.q2 ;
 wire \u_ro_only.ro_gen[2].ro2.q3 ;
 wire \u_ro_only.ro_gen[2].ro2.q4 ;
 wire \u_ro_only.ro_gen[3].ro1.cq4 ;
 wire \u_ro_only.ro_gen[3].ro1.q ;
 wire \u_ro_only.ro_gen[3].ro1.q0 ;
 wire \u_ro_only.ro_gen[3].ro1.q1 ;
 wire \u_ro_only.ro_gen[3].ro1.q2 ;
 wire \u_ro_only.ro_gen[3].ro1.q3 ;
 wire \u_ro_only.ro_gen[3].ro1.q4 ;
 wire \u_ro_only.ro_gen[3].ro2.cq4 ;
 wire \u_ro_only.ro_gen[3].ro2.q ;
 wire \u_ro_only.ro_gen[3].ro2.q0 ;
 wire \u_ro_only.ro_gen[3].ro2.q1 ;
 wire \u_ro_only.ro_gen[3].ro2.q2 ;
 wire \u_ro_only.ro_gen[3].ro2.q3 ;
 wire \u_ro_only.ro_gen[3].ro2.q4 ;
 wire \u_ro_only.ro_gen[4].ro1.cq4 ;
 wire \u_ro_only.ro_gen[4].ro1.q ;
 wire \u_ro_only.ro_gen[4].ro1.q0 ;
 wire \u_ro_only.ro_gen[4].ro1.q1 ;
 wire \u_ro_only.ro_gen[4].ro1.q2 ;
 wire \u_ro_only.ro_gen[4].ro1.q3 ;
 wire \u_ro_only.ro_gen[4].ro1.q4 ;
 wire \u_ro_only.ro_gen[4].ro2.cq4 ;
 wire \u_ro_only.ro_gen[4].ro2.q ;
 wire \u_ro_only.ro_gen[4].ro2.q0 ;
 wire \u_ro_only.ro_gen[4].ro2.q1 ;
 wire \u_ro_only.ro_gen[4].ro2.q2 ;
 wire \u_ro_only.ro_gen[4].ro2.q3 ;
 wire \u_ro_only.ro_gen[4].ro2.q4 ;
 wire \u_ro_only.ro_gen[5].ro1.cq4 ;
 wire \u_ro_only.ro_gen[5].ro1.q ;
 wire \u_ro_only.ro_gen[5].ro1.q0 ;
 wire \u_ro_only.ro_gen[5].ro1.q1 ;
 wire \u_ro_only.ro_gen[5].ro1.q2 ;
 wire \u_ro_only.ro_gen[5].ro1.q3 ;
 wire \u_ro_only.ro_gen[5].ro1.q4 ;
 wire \u_ro_only.ro_gen[5].ro2.cq4 ;
 wire \u_ro_only.ro_gen[5].ro2.q ;
 wire \u_ro_only.ro_gen[5].ro2.q0 ;
 wire \u_ro_only.ro_gen[5].ro2.q1 ;
 wire \u_ro_only.ro_gen[5].ro2.q2 ;
 wire \u_ro_only.ro_gen[5].ro2.q3 ;
 wire \u_ro_only.ro_gen[5].ro2.q4 ;
 wire \u_ro_only.ro_gen[6].ro1.cq4 ;
 wire \u_ro_only.ro_gen[6].ro1.q ;
 wire \u_ro_only.ro_gen[6].ro1.q0 ;
 wire \u_ro_only.ro_gen[6].ro1.q1 ;
 wire \u_ro_only.ro_gen[6].ro1.q2 ;
 wire \u_ro_only.ro_gen[6].ro1.q3 ;
 wire \u_ro_only.ro_gen[6].ro1.q4 ;
 wire \u_ro_only.ro_gen[6].ro2.cq4 ;
 wire \u_ro_only.ro_gen[6].ro2.q ;
 wire \u_ro_only.ro_gen[6].ro2.q0 ;
 wire \u_ro_only.ro_gen[6].ro2.q1 ;
 wire \u_ro_only.ro_gen[6].ro2.q2 ;
 wire \u_ro_only.ro_gen[6].ro2.q3 ;
 wire \u_ro_only.ro_gen[6].ro2.q4 ;
 wire \u_ro_only.ro_gen[7].ro1.cq4 ;
 wire \u_ro_only.ro_gen[7].ro1.q ;
 wire \u_ro_only.ro_gen[7].ro1.q0 ;
 wire \u_ro_only.ro_gen[7].ro1.q1 ;
 wire \u_ro_only.ro_gen[7].ro1.q2 ;
 wire \u_ro_only.ro_gen[7].ro1.q3 ;
 wire \u_ro_only.ro_gen[7].ro1.q4 ;
 wire \u_ro_only.ro_gen[7].ro2.cq4 ;
 wire \u_ro_only.ro_gen[7].ro2.q ;
 wire \u_ro_only.ro_gen[7].ro2.q0 ;
 wire \u_ro_only.ro_gen[7].ro2.q1 ;
 wire \u_ro_only.ro_gen[7].ro2.q2 ;
 wire \u_ro_only.ro_gen[7].ro2.q3 ;
 wire \u_ro_only.ro_gen[7].ro2.q4 ;
 wire \u_ro_only.ro_gen[8].ro1.cq4 ;
 wire \u_ro_only.ro_gen[8].ro1.q ;
 wire \u_ro_only.ro_gen[8].ro1.q0 ;
 wire \u_ro_only.ro_gen[8].ro1.q1 ;
 wire \u_ro_only.ro_gen[8].ro1.q2 ;
 wire \u_ro_only.ro_gen[8].ro1.q3 ;
 wire \u_ro_only.ro_gen[8].ro1.q4 ;
 wire \u_ro_only.ro_gen[8].ro2.cq4 ;
 wire \u_ro_only.ro_gen[8].ro2.q ;
 wire \u_ro_only.ro_gen[8].ro2.q0 ;
 wire \u_ro_only.ro_gen[8].ro2.q1 ;
 wire \u_ro_only.ro_gen[8].ro2.q2 ;
 wire \u_ro_only.ro_gen[8].ro2.q3 ;
 wire \u_ro_only.ro_gen[8].ro2.q4 ;
 wire \u_ro_only.ro_gen[9].ro1.cq4 ;
 wire \u_ro_only.ro_gen[9].ro1.q ;
 wire \u_ro_only.ro_gen[9].ro1.q0 ;
 wire \u_ro_only.ro_gen[9].ro1.q1 ;
 wire \u_ro_only.ro_gen[9].ro1.q2 ;
 wire \u_ro_only.ro_gen[9].ro1.q3 ;
 wire \u_ro_only.ro_gen[9].ro1.q4 ;
 wire \u_ro_only.ro_gen[9].ro2.cq4 ;
 wire \u_ro_only.ro_gen[9].ro2.q ;
 wire \u_ro_only.ro_gen[9].ro2.q0 ;
 wire \u_ro_only.ro_gen[9].ro2.q1 ;
 wire \u_ro_only.ro_gen[9].ro2.q2 ;
 wire \u_ro_only.ro_gen[9].ro2.q3 ;
 wire \u_ro_only.ro_gen[9].ro2.q4 ;
 wire clknet_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 sky130_fd_sc_hd__inv_2 _02_ (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00_));
 sky130_fd_sc_hd__and2_1 _03_ (.A(\u_ro_only.ro_gen[9].ro2.q ),
    .B(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[9].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _04_ (.A(\u_ro_only.ro_gen[9].ro1.q ),
    .B(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[9].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _05_ (.A(net6),
    .B(\u_ro_only.ro_gen[8].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[8].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _06_ (.A(net4),
    .B(\u_ro_only.ro_gen[8].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[8].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _07_ (.A(net7),
    .B(\u_ro_only.ro_gen[7].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[7].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _08_ (.A(net4),
    .B(\u_ro_only.ro_gen[7].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[7].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _09_ (.A(net6),
    .B(\u_ro_only.ro_gen[6].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[6].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _10_ (.A(net4),
    .B(\u_ro_only.ro_gen[6].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[6].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _11_ (.A(net6),
    .B(\u_ro_only.ro_gen[5].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[5].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _12_ (.A(net5),
    .B(\u_ro_only.ro_gen[5].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[5].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _13_ (.A(net7),
    .B(\u_ro_only.ro_gen[4].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[4].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _14_ (.A(net5),
    .B(\u_ro_only.ro_gen[4].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[4].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _15_ (.A(net6),
    .B(\u_ro_only.ro_gen[3].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[3].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _16_ (.A(net4),
    .B(\u_ro_only.ro_gen[3].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[3].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _17_ (.A(net6),
    .B(\u_ro_only.ro_gen[2].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[2].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _18_ (.A(net4),
    .B(\u_ro_only.ro_gen[2].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[2].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _19_ (.A(net7),
    .B(\u_ro_only.ro_gen[1].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[1].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _20_ (.A(net5),
    .B(\u_ro_only.ro_gen[1].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[1].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _21_ (.A(net6),
    .B(\u_ro_only.ro_gen[0].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[0].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _22_ (.A(net4),
    .B(\u_ro_only.ro_gen[0].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[0].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _23_ (.A(net7),
    .B(\u_ro_only.ro_gen[15].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[15].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _24_ (.A(net5),
    .B(\u_ro_only.ro_gen[15].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[15].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _25_ (.A(net6),
    .B(\u_ro_only.ro_gen[14].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[14].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _26_ (.A(net5),
    .B(\u_ro_only.ro_gen[14].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[14].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _27_ (.A(net6),
    .B(\u_ro_only.ro_gen[13].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[13].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _28_ (.A(net4),
    .B(\u_ro_only.ro_gen[13].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[13].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _29_ (.A(net6),
    .B(\u_ro_only.ro_gen[12].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[12].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _30_ (.A(net5),
    .B(\u_ro_only.ro_gen[12].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[12].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _31_ (.A(net7),
    .B(\u_ro_only.ro_gen[11].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[11].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _32_ (.A(net4),
    .B(\u_ro_only.ro_gen[11].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[11].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _33_ (.A(net7),
    .B(\u_ro_only.ro_gen[10].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[10].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _34_ (.A(net4),
    .B(\u_ro_only.ro_gen[10].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[10].ro1.cq4 ));
 sky130_fd_sc_hd__inv_2 _35_ (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01_));
 sky130_fd_sc_hd__dfrtp_1 _36_ (.CLK(clknet_1_1__leaf_clk),
    .D(net3),
    .RESET_B(_00_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_ro_only.ro_gen[0].ro2.en ));
 sky130_fd_sc_hd__dfrtp_1 _37_ (.CLK(clknet_1_0__leaf_clk),
    .D(net2),
    .RESET_B(_01_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_ro_only.ro_gen[0].ro1.en ));
 sky130_fd_sc_hd__buf_2 _38_ (.A(\u_ro_only.ro_gen[0].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[0].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _39_ (.A(\u_ro_only.ro_gen[0].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[0].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _40_ (.A(\u_ro_only.ro_gen[10].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[10].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _41_ (.A(\u_ro_only.ro_gen[10].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[10].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _42_ (.A(\u_ro_only.ro_gen[11].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[11].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _43_ (.A(\u_ro_only.ro_gen[11].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[11].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _44_ (.A(\u_ro_only.ro_gen[12].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[12].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _45_ (.A(\u_ro_only.ro_gen[12].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[12].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _46_ (.A(\u_ro_only.ro_gen[13].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[13].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _47_ (.A(\u_ro_only.ro_gen[13].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[13].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _48_ (.A(\u_ro_only.ro_gen[14].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[14].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _49_ (.A(\u_ro_only.ro_gen[14].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[14].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _50_ (.A(\u_ro_only.ro_gen[15].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[15].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _51_ (.A(\u_ro_only.ro_gen[15].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[15].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _52_ (.A(\u_ro_only.ro_gen[1].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[1].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _53_ (.A(\u_ro_only.ro_gen[1].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[1].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _54_ (.A(\u_ro_only.ro_gen[2].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[2].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _55_ (.A(\u_ro_only.ro_gen[2].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[2].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _56_ (.A(\u_ro_only.ro_gen[3].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[3].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _57_ (.A(\u_ro_only.ro_gen[3].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[3].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _58_ (.A(\u_ro_only.ro_gen[4].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[4].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _59_ (.A(\u_ro_only.ro_gen[4].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[4].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _60_ (.A(\u_ro_only.ro_gen[5].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[5].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _61_ (.A(\u_ro_only.ro_gen[5].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[5].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _62_ (.A(\u_ro_only.ro_gen[6].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[6].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _63_ (.A(\u_ro_only.ro_gen[6].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[6].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _64_ (.A(\u_ro_only.ro_gen[7].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[7].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _65_ (.A(\u_ro_only.ro_gen[7].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[7].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _66_ (.A(\u_ro_only.ro_gen[8].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[8].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _67_ (.A(\u_ro_only.ro_gen[8].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[8].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _68_ (.A(\u_ro_only.ro_gen[9].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[9].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _69_ (.A(\u_ro_only.ro_gen[9].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[9].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _70_ (.A(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[0]));
 sky130_fd_sc_hd__buf_2 _71_ (.A(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[1]));
 sky130_fd_sc_hd__buf_2 _72_ (.A(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[2]));
 sky130_fd_sc_hd__buf_2 _73_ (.A(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[3]));
 sky130_fd_sc_hd__buf_2 _74_ (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[4]));
 sky130_fd_sc_hd__buf_2 _75_ (.A(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[5]));
 sky130_fd_sc_hd__buf_2 _76_ (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[6]));
 sky130_fd_sc_hd__buf_2 _77_ (.A(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[7]));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[0].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[0].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[0].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[0].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[0].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[0].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[0].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[0].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[0].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[0].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[0].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[0].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[0].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[0].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[0].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[0].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[0].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[0].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[0].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[0].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[0].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[0].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[0].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[0].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[0].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[0].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[0].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[0].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[0].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[0].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[10].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[10].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[10].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[10].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[10].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[10].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[10].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[10].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[10].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[10].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[10].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[10].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[10].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[10].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[10].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[10].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[10].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[10].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[10].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[10].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[10].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[10].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[10].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[10].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[10].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[10].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[10].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[10].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[10].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[10].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[11].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[11].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[11].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[11].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[11].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[11].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[11].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[11].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[11].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[11].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[11].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[11].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[11].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[11].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[11].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[11].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[11].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[11].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[11].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[11].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[11].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[11].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[11].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[11].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[11].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[11].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[11].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[11].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[11].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[11].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[12].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[12].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[12].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[12].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[12].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[12].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[12].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[12].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[12].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[12].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[12].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[12].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[12].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[12].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[12].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[12].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[12].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[12].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[12].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[12].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[12].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[12].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[12].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[12].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[12].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[12].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[12].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[12].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[12].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[12].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[13].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[13].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[13].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[13].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[13].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[13].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[13].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[13].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[13].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[13].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[13].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[13].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[13].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[13].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[13].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[13].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[13].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[13].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[13].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[13].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[13].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[13].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[13].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[13].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[13].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[13].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[13].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[13].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[13].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[13].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[14].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[14].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[14].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[14].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[14].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[14].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[14].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[14].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[14].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[14].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[14].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[14].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[14].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[14].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[14].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[14].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[14].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[14].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[14].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[14].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[14].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[14].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[14].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[14].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[14].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[14].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[14].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[14].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[14].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[14].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[15].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[15].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[15].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[15].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[15].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[15].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[15].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[15].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[15].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[15].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[15].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[15].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[15].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[15].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[15].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[15].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[15].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[15].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[15].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[15].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[15].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[15].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[15].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[15].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[15].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[15].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[15].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[15].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[15].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[15].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[1].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[1].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[1].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[1].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[1].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[1].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[1].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[1].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[1].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[1].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[1].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[1].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[1].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[1].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[1].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[1].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[1].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[1].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[1].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[1].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[1].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[1].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[1].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[1].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[1].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[1].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[1].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[1].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[1].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[1].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[2].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[2].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[2].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[2].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[2].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[2].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[2].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[2].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[2].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[2].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[2].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[2].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[2].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[2].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[2].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[2].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[2].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[2].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[2].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[2].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[2].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[2].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[2].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[2].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[2].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[2].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[2].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[2].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[2].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[2].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[3].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[3].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[3].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[3].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[3].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[3].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[3].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[3].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[3].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[3].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[3].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[3].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[3].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[3].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[3].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[3].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[3].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[3].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[3].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[3].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[3].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[3].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[3].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[3].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[3].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[3].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[3].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[3].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[3].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[3].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[4].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[4].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[4].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[4].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[4].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[4].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[4].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[4].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[4].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[4].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[4].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[4].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[4].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[4].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[4].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[4].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[4].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[4].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[4].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[4].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[4].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[4].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[4].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[4].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[4].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[4].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[4].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[4].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[4].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[4].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[5].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[5].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[5].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[5].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[5].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[5].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[5].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[5].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[5].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[5].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[5].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[5].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[5].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[5].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[5].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[5].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[5].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[5].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[5].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[5].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[5].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[5].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[5].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[5].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[5].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[5].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[5].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[5].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[5].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[5].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[6].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[6].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[6].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[6].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[6].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[6].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[6].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[6].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[6].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[6].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[6].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[6].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[6].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[6].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[6].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[6].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[6].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[6].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[6].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[6].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[6].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[6].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[6].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[6].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[6].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[6].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[6].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[6].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[6].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[6].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[7].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[7].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[7].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[7].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[7].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[7].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[7].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[7].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[7].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[7].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[7].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[7].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[7].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[7].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[7].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[7].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[7].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[7].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[7].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[7].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[7].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[7].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[7].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[7].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[7].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[7].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[7].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[7].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[7].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[7].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[8].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[8].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[8].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[8].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[8].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[8].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[8].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[8].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[8].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[8].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[8].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[8].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[8].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[8].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[8].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[8].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[8].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[8].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[8].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[8].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[8].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[8].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[8].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[8].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[8].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[8].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[8].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[8].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[8].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[8].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[9].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[9].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[9].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[9].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[9].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[9].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[9].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[9].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[9].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[9].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[9].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[9].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[9].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[9].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[9].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[9].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[9].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[9].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[9].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[9].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[9].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[9].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[9].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[9].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[9].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[9].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[9].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[9].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[9].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[9].ro2.q ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__buf_1 input1 (.A(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ui_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 fanout4 (.A(\u_ro_only.ro_gen[0].ro1.en ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__buf_1 fanout5 (.A(\u_ro_only.ro_gen[0].ro1.en ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 fanout6 (.A(\u_ro_only.ro_gen[0].ro2.en ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__buf_1 fanout7 (.A(\u_ro_only.ro_gen[0].ro2.en ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__conb_1 _70__8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net8));
 sky130_fd_sc_hd__conb_1 _71__9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net9));
 sky130_fd_sc_hd__conb_1 _72__10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net10));
 sky130_fd_sc_hd__conb_1 _73__11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net11));
 sky130_fd_sc_hd__conb_1 _74__12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net12));
 sky130_fd_sc_hd__conb_1 _75__13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net13));
 sky130_fd_sc_hd__conb_1 _76__14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net14));
 sky130_fd_sc_hd__conb_1 _77__15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net15));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_clk));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_32 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_48 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_60 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_59 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_68 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_90 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_102 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_64 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
endmodule
