module tt_um_roy1707018_ro2 (clk,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uo_out);
 input clk;
 input rst_n;
 input VPWR;
 input VGND;
 input [7:0] ui_in;
 output [7:0] uo_out;

 wire \u_ro_only.ro_gen[0].ro1.cq4 ;
 wire \u_ro_only.ro_gen[0].ro1.en ;
 wire \u_ro_only.ro_gen[0].ro1.q ;
 wire \u_ro_only.ro_gen[0].ro1.q0 ;
 wire \u_ro_only.ro_gen[0].ro1.q1 ;
 wire \u_ro_only.ro_gen[0].ro1.q2 ;
 wire \u_ro_only.ro_gen[0].ro1.q3 ;
 wire \u_ro_only.ro_gen[0].ro1.q4 ;
 wire \u_ro_only.ro_gen[0].ro2.cq4 ;
 wire \u_ro_only.ro_gen[0].ro2.en ;
 wire \u_ro_only.ro_gen[0].ro2.q ;
 wire \u_ro_only.ro_gen[0].ro2.q0 ;
 wire \u_ro_only.ro_gen[0].ro2.q1 ;
 wire \u_ro_only.ro_gen[0].ro2.q2 ;
 wire \u_ro_only.ro_gen[0].ro2.q3 ;
 wire \u_ro_only.ro_gen[0].ro2.q4 ;
 wire \u_ro_only.ro_gen[1].ro1.cq4 ;
 wire \u_ro_only.ro_gen[1].ro1.q ;
 wire \u_ro_only.ro_gen[1].ro1.q0 ;
 wire \u_ro_only.ro_gen[1].ro1.q1 ;
 wire \u_ro_only.ro_gen[1].ro1.q2 ;
 wire \u_ro_only.ro_gen[1].ro1.q3 ;
 wire \u_ro_only.ro_gen[1].ro1.q4 ;
 wire \u_ro_only.ro_gen[1].ro2.cq4 ;
 wire \u_ro_only.ro_gen[1].ro2.q ;
 wire \u_ro_only.ro_gen[1].ro2.q0 ;
 wire \u_ro_only.ro_gen[1].ro2.q1 ;
 wire \u_ro_only.ro_gen[1].ro2.q2 ;
 wire \u_ro_only.ro_gen[1].ro2.q3 ;
 wire \u_ro_only.ro_gen[1].ro2.q4 ;
 wire \u_ro_only.ro_gen[2].ro1.cq4 ;
 wire \u_ro_only.ro_gen[2].ro1.q ;
 wire \u_ro_only.ro_gen[2].ro1.q0 ;
 wire \u_ro_only.ro_gen[2].ro1.q1 ;
 wire \u_ro_only.ro_gen[2].ro1.q2 ;
 wire \u_ro_only.ro_gen[2].ro1.q3 ;
 wire \u_ro_only.ro_gen[2].ro1.q4 ;
 wire \u_ro_only.ro_gen[2].ro2.cq4 ;
 wire \u_ro_only.ro_gen[2].ro2.q ;
 wire \u_ro_only.ro_gen[2].ro2.q0 ;
 wire \u_ro_only.ro_gen[2].ro2.q1 ;
 wire \u_ro_only.ro_gen[2].ro2.q2 ;
 wire \u_ro_only.ro_gen[2].ro2.q3 ;
 wire \u_ro_only.ro_gen[2].ro2.q4 ;
 wire \u_ro_only.ro_gen[3].ro1.cq4 ;
 wire \u_ro_only.ro_gen[3].ro1.q ;
 wire \u_ro_only.ro_gen[3].ro1.q0 ;
 wire \u_ro_only.ro_gen[3].ro1.q1 ;
 wire \u_ro_only.ro_gen[3].ro1.q2 ;
 wire \u_ro_only.ro_gen[3].ro1.q3 ;
 wire \u_ro_only.ro_gen[3].ro1.q4 ;
 wire \u_ro_only.ro_gen[3].ro2.cq4 ;
 wire \u_ro_only.ro_gen[3].ro2.q ;
 wire \u_ro_only.ro_gen[3].ro2.q0 ;
 wire \u_ro_only.ro_gen[3].ro2.q1 ;
 wire \u_ro_only.ro_gen[3].ro2.q2 ;
 wire \u_ro_only.ro_gen[3].ro2.q3 ;
 wire \u_ro_only.ro_gen[3].ro2.q4 ;
 wire \u_ro_only.ro_gen[4].ro1.cq4 ;
 wire \u_ro_only.ro_gen[4].ro1.q ;
 wire \u_ro_only.ro_gen[4].ro1.q0 ;
 wire \u_ro_only.ro_gen[4].ro1.q1 ;
 wire \u_ro_only.ro_gen[4].ro1.q2 ;
 wire \u_ro_only.ro_gen[4].ro1.q3 ;
 wire \u_ro_only.ro_gen[4].ro1.q4 ;
 wire \u_ro_only.ro_gen[4].ro2.cq4 ;
 wire \u_ro_only.ro_gen[4].ro2.q ;
 wire \u_ro_only.ro_gen[4].ro2.q0 ;
 wire \u_ro_only.ro_gen[4].ro2.q1 ;
 wire \u_ro_only.ro_gen[4].ro2.q2 ;
 wire \u_ro_only.ro_gen[4].ro2.q3 ;
 wire \u_ro_only.ro_gen[4].ro2.q4 ;
 wire \u_ro_only.ro_gen[5].ro1.cq4 ;
 wire \u_ro_only.ro_gen[5].ro1.q ;
 wire \u_ro_only.ro_gen[5].ro1.q0 ;
 wire \u_ro_only.ro_gen[5].ro1.q1 ;
 wire \u_ro_only.ro_gen[5].ro1.q2 ;
 wire \u_ro_only.ro_gen[5].ro1.q3 ;
 wire \u_ro_only.ro_gen[5].ro1.q4 ;
 wire \u_ro_only.ro_gen[5].ro2.cq4 ;
 wire \u_ro_only.ro_gen[5].ro2.q ;
 wire \u_ro_only.ro_gen[5].ro2.q0 ;
 wire \u_ro_only.ro_gen[5].ro2.q1 ;
 wire \u_ro_only.ro_gen[5].ro2.q2 ;
 wire \u_ro_only.ro_gen[5].ro2.q3 ;
 wire \u_ro_only.ro_gen[5].ro2.q4 ;
 wire \u_ro_only.ro_gen[6].ro1.cq4 ;
 wire \u_ro_only.ro_gen[6].ro1.q ;
 wire \u_ro_only.ro_gen[6].ro1.q0 ;
 wire \u_ro_only.ro_gen[6].ro1.q1 ;
 wire \u_ro_only.ro_gen[6].ro1.q2 ;
 wire \u_ro_only.ro_gen[6].ro1.q3 ;
 wire \u_ro_only.ro_gen[6].ro1.q4 ;
 wire \u_ro_only.ro_gen[6].ro2.cq4 ;
 wire \u_ro_only.ro_gen[6].ro2.q ;
 wire \u_ro_only.ro_gen[6].ro2.q0 ;
 wire \u_ro_only.ro_gen[6].ro2.q1 ;
 wire \u_ro_only.ro_gen[6].ro2.q2 ;
 wire \u_ro_only.ro_gen[6].ro2.q3 ;
 wire \u_ro_only.ro_gen[6].ro2.q4 ;
 wire \u_ro_only.ro_gen[7].ro1.cq4 ;
 wire \u_ro_only.ro_gen[7].ro1.q ;
 wire \u_ro_only.ro_gen[7].ro1.q0 ;
 wire \u_ro_only.ro_gen[7].ro1.q1 ;
 wire \u_ro_only.ro_gen[7].ro1.q2 ;
 wire \u_ro_only.ro_gen[7].ro1.q3 ;
 wire \u_ro_only.ro_gen[7].ro1.q4 ;
 wire \u_ro_only.ro_gen[7].ro2.cq4 ;
 wire \u_ro_only.ro_gen[7].ro2.q ;
 wire \u_ro_only.ro_gen[7].ro2.q0 ;
 wire \u_ro_only.ro_gen[7].ro2.q1 ;
 wire \u_ro_only.ro_gen[7].ro2.q2 ;
 wire \u_ro_only.ro_gen[7].ro2.q3 ;
 wire \u_ro_only.ro_gen[7].ro2.q4 ;
 wire clknet_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 sky130_fd_sc_hd__and2_1 _00_ (.A(\u_ro_only.ro_gen[1].ro1.q ),
    .B(\u_ro_only.ro_gen[0].ro1.en ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[1].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _01_ (.A(\u_ro_only.ro_gen[0].ro2.q ),
    .B(\u_ro_only.ro_gen[0].ro2.en ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[0].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _02_ (.A(\u_ro_only.ro_gen[0].ro1.en ),
    .B(\u_ro_only.ro_gen[0].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[0].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _03_ (.A(\u_ro_only.ro_gen[0].ro2.en ),
    .B(\u_ro_only.ro_gen[7].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[7].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _04_ (.A(\u_ro_only.ro_gen[0].ro1.en ),
    .B(\u_ro_only.ro_gen[7].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[7].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _05_ (.A(\u_ro_only.ro_gen[0].ro2.en ),
    .B(\u_ro_only.ro_gen[6].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[6].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _06_ (.A(\u_ro_only.ro_gen[0].ro1.en ),
    .B(\u_ro_only.ro_gen[6].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[6].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _07_ (.A(\u_ro_only.ro_gen[0].ro2.en ),
    .B(\u_ro_only.ro_gen[5].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[5].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _08_ (.A(\u_ro_only.ro_gen[0].ro1.en ),
    .B(\u_ro_only.ro_gen[5].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[5].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _09_ (.A(\u_ro_only.ro_gen[0].ro2.en ),
    .B(\u_ro_only.ro_gen[4].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[4].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _10_ (.A(\u_ro_only.ro_gen[0].ro1.en ),
    .B(\u_ro_only.ro_gen[4].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[4].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _11_ (.A(\u_ro_only.ro_gen[0].ro2.en ),
    .B(\u_ro_only.ro_gen[3].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[3].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _12_ (.A(\u_ro_only.ro_gen[0].ro1.en ),
    .B(\u_ro_only.ro_gen[3].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[3].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _13_ (.A(\u_ro_only.ro_gen[0].ro2.en ),
    .B(\u_ro_only.ro_gen[2].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[2].ro2.cq4 ));
 sky130_fd_sc_hd__and2_1 _14_ (.A(\u_ro_only.ro_gen[0].ro1.en ),
    .B(\u_ro_only.ro_gen[2].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[2].ro1.cq4 ));
 sky130_fd_sc_hd__and2_1 _15_ (.A(\u_ro_only.ro_gen[0].ro2.en ),
    .B(\u_ro_only.ro_gen[1].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[1].ro2.cq4 ));
 sky130_fd_sc_hd__dfxtp_1 _16_ (.CLK(clknet_1_0__leaf_clk),
    .D(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_ro_only.ro_gen[0].ro1.en ));
 sky130_fd_sc_hd__dfxtp_1 _17_ (.CLK(clknet_1_1__leaf_clk),
    .D(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\u_ro_only.ro_gen[0].ro2.en ));
 sky130_fd_sc_hd__buf_2 _18_ (.A(\u_ro_only.ro_gen[0].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[0].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _19_ (.A(\u_ro_only.ro_gen[0].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[0].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _20_ (.A(\u_ro_only.ro_gen[1].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[1].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _21_ (.A(\u_ro_only.ro_gen[1].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[1].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _22_ (.A(\u_ro_only.ro_gen[2].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[2].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _23_ (.A(\u_ro_only.ro_gen[2].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[2].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _24_ (.A(\u_ro_only.ro_gen[3].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[3].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _25_ (.A(\u_ro_only.ro_gen[3].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[3].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _26_ (.A(\u_ro_only.ro_gen[4].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[4].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _27_ (.A(\u_ro_only.ro_gen[4].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[4].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _28_ (.A(\u_ro_only.ro_gen[5].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[5].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _29_ (.A(\u_ro_only.ro_gen[5].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[5].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _30_ (.A(\u_ro_only.ro_gen[6].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[6].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _31_ (.A(\u_ro_only.ro_gen[6].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[6].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _32_ (.A(\u_ro_only.ro_gen[7].ro1.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[7].ro1.q4 ));
 sky130_fd_sc_hd__buf_2 _33_ (.A(\u_ro_only.ro_gen[7].ro2.q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\u_ro_only.ro_gen[7].ro2.q4 ));
 sky130_fd_sc_hd__buf_2 _34_ (.A(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[0]));
 sky130_fd_sc_hd__buf_2 _35_ (.A(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[1]));
 sky130_fd_sc_hd__buf_2 _36_ (.A(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[2]));
 sky130_fd_sc_hd__buf_2 _37_ (.A(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[3]));
 sky130_fd_sc_hd__buf_2 _38_ (.A(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[4]));
 sky130_fd_sc_hd__buf_2 _39_ (.A(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[5]));
 sky130_fd_sc_hd__buf_2 _40_ (.A(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[6]));
 sky130_fd_sc_hd__buf_2 _41_ (.A(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[7]));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[0].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[0].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[0].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[0].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[0].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[0].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[0].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[0].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[0].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[0].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[0].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[0].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[0].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[0].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[0].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[0].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[0].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[0].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[0].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[0].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[0].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[0].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[0].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[0].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[0].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[0].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[0].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[0].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[0].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[0].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[1].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[1].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[1].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[1].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[1].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[1].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[1].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[1].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[1].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[1].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[1].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[1].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[1].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[1].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[1].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[1].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[1].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[1].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[1].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[1].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[1].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[1].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[1].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[1].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[1].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[1].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[1].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[1].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[1].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[1].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[2].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[2].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[2].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[2].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[2].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[2].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[2].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[2].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[2].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[2].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[2].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[2].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[2].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[2].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[2].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[2].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[2].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[2].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[2].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[2].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[2].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[2].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[2].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[2].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[2].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[2].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[2].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[2].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[2].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[2].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[3].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[3].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[3].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[3].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[3].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[3].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[3].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[3].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[3].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[3].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[3].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[3].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[3].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[3].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[3].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[3].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[3].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[3].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[3].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[3].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[3].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[3].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[3].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[3].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[3].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[3].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[3].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[3].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[3].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[3].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[4].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[4].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[4].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[4].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[4].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[4].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[4].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[4].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[4].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[4].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[4].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[4].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[4].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[4].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[4].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[4].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[4].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[4].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[4].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[4].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[4].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[4].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[4].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[4].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[4].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[4].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[4].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[4].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[4].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[4].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[5].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[5].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[5].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[5].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[5].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[5].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[5].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[5].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[5].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[5].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[5].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[5].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[5].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[5].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[5].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[5].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[5].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[5].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[5].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[5].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[5].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[5].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[5].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[5].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[5].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[5].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[5].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[5].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[5].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[5].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[6].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[6].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[6].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[6].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[6].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[6].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[6].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[6].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[6].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[6].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[6].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[6].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[6].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[6].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[6].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[6].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[6].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[6].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[6].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[6].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[6].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[6].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[6].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[6].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[6].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[6].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[6].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[6].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[6].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[6].ro2.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[7].ro1.cinv1/_0_  (.A(\u_ro_only.ro_gen[7].ro1.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[7].ro1.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[7].ro1.cinv2/_0_  (.A(\u_ro_only.ro_gen[7].ro1.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[7].ro1.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[7].ro1.cinv3/_0_  (.A(\u_ro_only.ro_gen[7].ro1.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[7].ro1.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[7].ro1.cinv4/_0_  (.A(\u_ro_only.ro_gen[7].ro1.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[7].ro1.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[7].ro1.cinv5/_0_  (.A(\u_ro_only.ro_gen[7].ro1.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[7].ro1.q ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[7].ro2.cinv1/_0_  (.A(\u_ro_only.ro_gen[7].ro2.cq4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[7].ro2.q0 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[7].ro2.cinv2/_0_  (.A(\u_ro_only.ro_gen[7].ro2.q0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[7].ro2.q1 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[7].ro2.cinv3/_0_  (.A(\u_ro_only.ro_gen[7].ro2.q1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[7].ro2.q2 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[7].ro2.cinv4/_0_  (.A(\u_ro_only.ro_gen[7].ro2.q2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[7].ro2.q3 ));
 sky130_fd_sc_hd__inv_2 \u_ro_only.ro_gen[7].ro2.cinv5/_0_  (.A(\u_ro_only.ro_gen[7].ro2.q3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\u_ro_only.ro_gen[7].ro2.q ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ui_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__conb_1 _34__3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net3));
 sky130_fd_sc_hd__conb_1 _35__4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net4));
 sky130_fd_sc_hd__conb_1 _36__5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net5));
 sky130_fd_sc_hd__conb_1 _37__6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net6));
 sky130_fd_sc_hd__conb_1 _38__7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net7));
 sky130_fd_sc_hd__conb_1 _39__8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net8));
 sky130_fd_sc_hd__conb_1 _40__9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net9));
 sky130_fd_sc_hd__conb_1 _41__10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net10));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_clk));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_44 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_91 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_91 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
endmodule
